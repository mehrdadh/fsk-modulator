/* Verilog model created from schematic test.sch -- May 22, 2019 17:58 */

module test;




endmodule // test
