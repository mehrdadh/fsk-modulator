/* Verilog model created from schematic test.sch -- May 22, 2019 13:46 */

module test;




endmodule // test
