module ble_mem(
	addr,
	data
);

input [7:0]	addr;
output reg	data;


endmodule