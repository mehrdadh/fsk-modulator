module ble_packet(addr, data);
input [9:0] addr;
output reg	[25:0] data;

reg [25:0] sineTable[0:1023];
always @(addr)
	data	=	sineTable[addr];

always begin
	sineTable[10'd0] = 26'b01111111111110000000000000;
	sineTable[10'd1] = 26'b01100100001000100111110101;
	sineTable[10'd2] = 26'b00000000000000111111111111;
	sineTable[10'd3] = 26'b10011011110110100111110101;
	sineTable[10'd4] = 26'b10000000000010000000000000;
	sineTable[10'd5] = 26'b10011011110110100111110101;
	sineTable[10'd6] = 26'b00000000000000111111111111;
	sineTable[10'd7] = 26'b01100100001000100111110101;
	sineTable[10'd8] = 26'b01111111111110000000000000;
	sineTable[10'd9] = 26'b01100100001000100111110101;
	sineTable[10'd10] = 26'b00000000000000111111111111;
	sineTable[10'd11] = 26'b10011011110110100111110101;
	sineTable[10'd12] = 26'b10000000000010000000000000;
	sineTable[10'd13] = 26'b10011011110110100111110101;
	sineTable[10'd14] = 26'b00000000000000111111111111;
	sineTable[10'd15] = 26'b01100100001000100111110101;
	sineTable[10'd16] = 26'b01111111111110000000000000;
	sineTable[10'd17] = 26'b01100100001000100111110101;
	sineTable[10'd18] = 26'b00000000000000111111111111;
	sineTable[10'd19] = 26'b10011011110110100111110101;
	sineTable[10'd20] = 26'b10000000000010000000000000;
	sineTable[10'd21] = 26'b10011011110110100111110101;
	sineTable[10'd22] = 26'b00000000000000111111111111;
	sineTable[10'd23] = 26'b01100100001000100111110101;
	sineTable[10'd24] = 26'b01111111111110000000000000;
	sineTable[10'd25] = 26'b01100100001000100111110101;
	sineTable[10'd26] = 26'b00000000000000111111111111;
	sineTable[10'd27] = 26'b10011011110110100111110101;
	sineTable[10'd28] = 26'b10000000000010000000000000;
	sineTable[10'd29] = 26'b10011011110110100111110101;
	sineTable[10'd30] = 26'b00000000000000111111111111;
	sineTable[10'd31] = 26'b01100100001000100111110101;
	sineTable[10'd32] = 26'b01111111111110000000000000;
	sineTable[10'd33] = 26'b01100100001000100111110101;
	sineTable[10'd34] = 26'b00000000000000111111111111;
	sineTable[10'd35] = 26'b10011011110110100111110101;
	sineTable[10'd36] = 26'b10000000000010000000000000;
	sineTable[10'd37] = 26'b10011011110110100111110101;
	sineTable[10'd38] = 26'b00000000000000111111111111;
	sineTable[10'd39] = 26'b01100100001000100111110101;
	sineTable[10'd40] = 26'b01111111111110000000000000;
	sineTable[10'd41] = 26'b01100100001001011000001010;
	sineTable[10'd42] = 26'b00000000000001000000000001;
	sineTable[10'd43] = 26'b10011011110111011000001010;
	sineTable[10'd44] = 26'b10000000000011111111111111;
	sineTable[10'd45] = 26'b10011011110111011000001010;
	sineTable[10'd46] = 26'b00000000000001000000000001;
	sineTable[10'd47] = 26'b01100100001001011000001010;
	sineTable[10'd48] = 26'b01111111111110000000000000;
	sineTable[10'd49] = 26'b01100100001001011000001010;
	sineTable[10'd50] = 26'b00000000000001000000000001;
	sineTable[10'd51] = 26'b10011011110111011000001010;
	sineTable[10'd52] = 26'b10000000000011111111111111;
	sineTable[10'd53] = 26'b10011011110111011000001010;
	sineTable[10'd54] = 26'b00000000000001000000000001;
	sineTable[10'd55] = 26'b01100100001001011000001010;
	sineTable[10'd56] = 26'b01111111111110000000000000;
	sineTable[10'd57] = 26'b01100100001001011000001010;
	sineTable[10'd58] = 26'b00000000000001000000000001;
	sineTable[10'd59] = 26'b10011011110111011000001010;
	sineTable[10'd60] = 26'b10000000000011111111111111;
	sineTable[10'd61] = 26'b10011011110110100111110101;
	sineTable[10'd62] = 26'b11111111111110111111111111;
	sineTable[10'd63] = 26'b01100100001000100111110101;
	sineTable[10'd64] = 26'b01111111111110000000000000;
	sineTable[10'd65] = 26'b01100100001000100111110101;
	sineTable[10'd66] = 26'b11111111111110111111111111;
	sineTable[10'd67] = 26'b10011011110110100111110101;
	sineTable[10'd68] = 26'b10000000000011111111111111;
	sineTable[10'd69] = 26'b10011011110110100111110101;
	sineTable[10'd70] = 26'b11111111111110111111111111;
	sineTable[10'd71] = 26'b01100100001000100111110101;
	sineTable[10'd72] = 26'b01111111111110000000000000;
	sineTable[10'd73] = 26'b01100100001001011000001010;
	sineTable[10'd74] = 26'b00000000000001000000000001;
	sineTable[10'd75] = 26'b10011011110111011000001010;
	sineTable[10'd76] = 26'b10000000000011111111111111;
	sineTable[10'd77] = 26'b10011011110110100111110101;
	sineTable[10'd78] = 26'b11111111111110111111111111;
	sineTable[10'd79] = 26'b01100100001000100111110101;
	sineTable[10'd80] = 26'b01111111111110000000000000;
	sineTable[10'd81] = 26'b01100100001001011000001010;
	sineTable[10'd82] = 26'b00000000000001000000000001;
	sineTable[10'd83] = 26'b10011011110111011000001010;
	sineTable[10'd84] = 26'b10000000000011111111111111;
	sineTable[10'd85] = 26'b10011011110110100111110101;
	sineTable[10'd86] = 26'b11111111111110111111111111;
	sineTable[10'd87] = 26'b01100100001000100111110101;
	sineTable[10'd88] = 26'b01111111111110000000000000;
	sineTable[10'd89] = 26'b01100100001000100111110101;
	sineTable[10'd90] = 26'b11111111111110111111111111;
	sineTable[10'd91] = 26'b10011011110110100111110101;
	sineTable[10'd92] = 26'b10000000000011111111111111;
	sineTable[10'd93] = 26'b10011011110110100111110101;
	sineTable[10'd94] = 26'b11111111111110111111111111;
	sineTable[10'd95] = 26'b01100100001000100111110101;
	sineTable[10'd96] = 26'b01111111111110000000000000;
	sineTable[10'd97] = 26'b01100100001001011000001010;
	sineTable[10'd98] = 26'b00000000000001000000000001;
	sineTable[10'd99] = 26'b10011011110111011000001010;
	sineTable[10'd100] = 26'b10000000000011111111111111;
	sineTable[10'd101] = 26'b10011011110111011000001010;
	sineTable[10'd102] = 26'b00000000000001000000000001;
	sineTable[10'd103] = 26'b01100100001001011000001010;
	sineTable[10'd104] = 26'b01111111111110000000000000;
	sineTable[10'd105] = 26'b01100100001000100111110101;
	sineTable[10'd106] = 26'b11111111111110111111111111;
	sineTable[10'd107] = 26'b10011011110110100111110101;
	sineTable[10'd108] = 26'b10000000000011111111111111;
	sineTable[10'd109] = 26'b10011011110110100111110101;
	sineTable[10'd110] = 26'b11111111111110111111111111;
	sineTable[10'd111] = 26'b01100100001000100111110101;
	sineTable[10'd112] = 26'b01111111111110000000000000;
	sineTable[10'd113] = 26'b01100100001000100111110101;
	sineTable[10'd114] = 26'b11111111111110111111111111;
	sineTable[10'd115] = 26'b10011011110110100111110101;
	sineTable[10'd116] = 26'b10000000000011111111111111;
	sineTable[10'd117] = 26'b10011011110111011000001010;
	sineTable[10'd118] = 26'b00000000000001000000000001;
	sineTable[10'd119] = 26'b01100100001001011000001010;
	sineTable[10'd120] = 26'b01111111111110000000000000;
	sineTable[10'd121] = 26'b01100100001000100111110101;
	sineTable[10'd122] = 26'b11111111111110111111111111;
	sineTable[10'd123] = 26'b10011011110110100111110101;
	sineTable[10'd124] = 26'b10000000000011111111111111;
	sineTable[10'd125] = 26'b10011011110110100111110101;
	sineTable[10'd126] = 26'b11111111111110111111111111;
	sineTable[10'd127] = 26'b01100100001000100111110101;
	sineTable[10'd128] = 26'b01111111111110000000000000;
	sineTable[10'd129] = 26'b01100100001000100111110101;
	sineTable[10'd130] = 26'b11111111111110111111111111;
	sineTable[10'd131] = 26'b10011011110110100111110101;
	sineTable[10'd132] = 26'b10000000000011111111111111;
	sineTable[10'd133] = 26'b10011011110110100111110101;
	sineTable[10'd134] = 26'b11111111111110111111111111;
	sineTable[10'd135] = 26'b01100100001000100111110101;
	sineTable[10'd136] = 26'b01111111111110000000000000;
	sineTable[10'd137] = 26'b01100100001001011000001010;
	sineTable[10'd138] = 26'b00000000000001000000000001;
	sineTable[10'd139] = 26'b10011011110111011000001010;
	sineTable[10'd140] = 26'b10000000000011111111111111;
	sineTable[10'd141] = 26'b10011011110110100111110101;
	sineTable[10'd142] = 26'b11111111111110111111111111;
	sineTable[10'd143] = 26'b01100100001000100111110101;
	sineTable[10'd144] = 26'b01111111111110000000000000;
	sineTable[10'd145] = 26'b01100100001000100111110101;
	sineTable[10'd146] = 26'b11111111111110111111111111;
	sineTable[10'd147] = 26'b10011011110110100111110101;
	sineTable[10'd148] = 26'b10000000000011111111111111;
	sineTable[10'd149] = 26'b10011011110111011000001010;
	sineTable[10'd150] = 26'b00000000000001000000000001;
	sineTable[10'd151] = 26'b01100100001001011000001010;
	sineTable[10'd152] = 26'b01111111111110000000000000;
	sineTable[10'd153] = 26'b01100100001000100111110101;
	sineTable[10'd154] = 26'b11111111111110111111111111;
	sineTable[10'd155] = 26'b10011011110110100111110101;
	sineTable[10'd156] = 26'b10000000000011111111111111;
	sineTable[10'd157] = 26'b10011011110110100111110101;
	sineTable[10'd158] = 26'b11111111111110111111111111;
	sineTable[10'd159] = 26'b01100100001000100111110101;
	sineTable[10'd160] = 26'b01111111111110000000000000;
	sineTable[10'd161] = 26'b01100100001000100111110101;
	sineTable[10'd162] = 26'b11111111111110111111111111;
	sineTable[10'd163] = 26'b10011011110110100111110101;
	sineTable[10'd164] = 26'b10000000000011111111111111;
	sineTable[10'd165] = 26'b10011011110110100111110101;
	sineTable[10'd166] = 26'b11111111111110111111111111;
	sineTable[10'd167] = 26'b01100100001000100111110101;
	sineTable[10'd168] = 26'b01111111111110000000000000;
	sineTable[10'd169] = 26'b01100100001001011000001010;
	sineTable[10'd170] = 26'b00000000000001000000000001;
	sineTable[10'd171] = 26'b10011011110111011000001010;
	sineTable[10'd172] = 26'b10000000000011111111111111;
	sineTable[10'd173] = 26'b10011011110111011000001010;
	sineTable[10'd174] = 26'b00000000000001000000000001;
	sineTable[10'd175] = 26'b01100100001001011000001010;
	sineTable[10'd176] = 26'b01111111111110000000000000;
	sineTable[10'd177] = 26'b01100100001000100111110101;
	sineTable[10'd178] = 26'b11111111111110111111111111;
	sineTable[10'd179] = 26'b10011011110110100111110101;
	sineTable[10'd180] = 26'b10000000000011111111111111;
	sineTable[10'd181] = 26'b10011011110111011000001010;
	sineTable[10'd182] = 26'b00000000000001000000000001;
	sineTable[10'd183] = 26'b01100100001001011000001010;
	sineTable[10'd184] = 26'b01111111111110000000000000;
	sineTable[10'd185] = 26'b01100100001001011000001010;
	sineTable[10'd186] = 26'b00000000000001000000000001;
	sineTable[10'd187] = 26'b10011011110111011000001010;
	sineTable[10'd188] = 26'b10000000000011111111111111;
	sineTable[10'd189] = 26'b10011011110111011000001010;
	sineTable[10'd190] = 26'b00000000000001000000000001;
	sineTable[10'd191] = 26'b01100100001001011000001010;
	sineTable[10'd192] = 26'b01111111111110000000000000;
	sineTable[10'd193] = 26'b01100100001000100111110101;
	sineTable[10'd194] = 26'b11111111111110111111111111;
	sineTable[10'd195] = 26'b10011011110110100111110101;
	sineTable[10'd196] = 26'b10000000000011111111111111;
	sineTable[10'd197] = 26'b10011011110110100111110101;
	sineTable[10'd198] = 26'b11111111111110111111111111;
	sineTable[10'd199] = 26'b01100100001000100111110101;
	sineTable[10'd200] = 26'b01111111111110000000000000;
	sineTable[10'd201] = 26'b01100100001001011000001010;
	sineTable[10'd202] = 26'b00000000000001000000000001;
	sineTable[10'd203] = 26'b10011011110111011000001010;
	sineTable[10'd204] = 26'b10000000000011111111111111;
	sineTable[10'd205] = 26'b10011011110111011000001010;
	sineTable[10'd206] = 26'b00000000000001000000000001;
	sineTable[10'd207] = 26'b01100100001001011000001010;
	sineTable[10'd208] = 26'b01111111111110000000000000;
	sineTable[10'd209] = 26'b01100100001001011000001010;
	sineTable[10'd210] = 26'b00000000000001000000000001;
	sineTable[10'd211] = 26'b10011011110111011000001010;
	sineTable[10'd212] = 26'b10000000000011111111111111;
	sineTable[10'd213] = 26'b10011011110110100111110101;
	sineTable[10'd214] = 26'b11111111111110111111111111;
	sineTable[10'd215] = 26'b01100100001000100111110101;
	sineTable[10'd216] = 26'b01111111111110000000000000;
	sineTable[10'd217] = 26'b01100100001000100111110101;
	sineTable[10'd218] = 26'b11111111111110111111111111;
	sineTable[10'd219] = 26'b10011011110110100111110101;
	sineTable[10'd220] = 26'b10000000000011111111111111;
	sineTable[10'd221] = 26'b10011011110111011000001010;
	sineTable[10'd222] = 26'b00000000000001000000000001;
	sineTable[10'd223] = 26'b01100100001001011000001010;
	sineTable[10'd224] = 26'b01111111111110000000000000;
	sineTable[10'd225] = 26'b01100100001000100111110101;
	sineTable[10'd226] = 26'b11111111111110111111111111;
	sineTable[10'd227] = 26'b10011011110110100111110101;
	sineTable[10'd228] = 26'b10000000000011111111111111;
	sineTable[10'd229] = 26'b10011011110111011000001010;
	sineTable[10'd230] = 26'b00000000000001000000000001;
	sineTable[10'd231] = 26'b01100100001001011000001010;
	sineTable[10'd232] = 26'b01111111111110000000000000;
	sineTable[10'd233] = 26'b01100100001000100111110101;
	sineTable[10'd234] = 26'b11111111111110111111111111;
	sineTable[10'd235] = 26'b10011011110110100111110101;
	sineTable[10'd236] = 26'b10000000000011111111111111;
	sineTable[10'd237] = 26'b10011011110110100111110101;
	sineTable[10'd238] = 26'b11111111111110111111111111;
	sineTable[10'd239] = 26'b01100100001000100111110101;
	sineTable[10'd240] = 26'b01111111111110000000000000;
	sineTable[10'd241] = 26'b01100100001001011000001010;
	sineTable[10'd242] = 26'b00000000000001000000000001;
	sineTable[10'd243] = 26'b10011011110111011000001010;
	sineTable[10'd244] = 26'b10000000000011111111111111;
	sineTable[10'd245] = 26'b10011011110111011000001010;
	sineTable[10'd246] = 26'b00000000000001000000000001;
	sineTable[10'd247] = 26'b01100100001001011000001010;
	sineTable[10'd248] = 26'b01111111111110000000000000;
	sineTable[10'd249] = 26'b01100100001001011000001010;
	sineTable[10'd250] = 26'b00000000000001000000000001;
	sineTable[10'd251] = 26'b10011011110111011000001010;
	sineTable[10'd252] = 26'b10000000000011111111111111;
	sineTable[10'd253] = 26'b10011011110111011000001010;
	sineTable[10'd254] = 26'b00000000000001000000000001;
	sineTable[10'd255] = 26'b01100100001001011000001010;
	sineTable[10'd256] = 26'b01111111111110000000000000;
	sineTable[10'd257] = 26'b01100100001000100111110101;
	sineTable[10'd258] = 26'b11111111111110111111111111;
	sineTable[10'd259] = 26'b10011011110110100111110101;
	sineTable[10'd260] = 26'b10000000000011111111111111;
	sineTable[10'd261] = 26'b10011011110111011000001010;
	sineTable[10'd262] = 26'b00000000000001000000000001;
	sineTable[10'd263] = 26'b01100100001001011000001010;
	sineTable[10'd264] = 26'b01111111111110000000000000;
	sineTable[10'd265] = 26'b01100100001001011000001010;
	sineTable[10'd266] = 26'b00000000000001000000000001;
	sineTable[10'd267] = 26'b10011011110111011000001010;
	sineTable[10'd268] = 26'b10000000000011111111111111;
	sineTable[10'd269] = 26'b10011011110110100111110101;
	sineTable[10'd270] = 26'b11111111111110111111111111;
	sineTable[10'd271] = 26'b01100100001000100111110101;
	sineTable[10'd272] = 26'b01111111111110000000000000;
	sineTable[10'd273] = 26'b01100100001001011000001010;
	sineTable[10'd274] = 26'b00000000000001000000000001;
	sineTable[10'd275] = 26'b10011011110111011000001010;
	sineTable[10'd276] = 26'b10000000000011111111111111;
	sineTable[10'd277] = 26'b10011011110111011000001010;
	sineTable[10'd278] = 26'b00000000000001000000000001;
	sineTable[10'd279] = 26'b01100100001001011000001010;
	sineTable[10'd280] = 26'b01111111111110000000000000;
	sineTable[10'd281] = 26'b01100100001001011000001010;
	sineTable[10'd282] = 26'b00000000000001000000000001;
	sineTable[10'd283] = 26'b10011011110111011000001010;
	sineTable[10'd284] = 26'b10000000000011111111111111;
	sineTable[10'd285] = 26'b10011011110110100111110101;
	sineTable[10'd286] = 26'b11111111111110111111111111;
	sineTable[10'd287] = 26'b01100100001000100111110101;
	sineTable[10'd288] = 26'b01111111111110000000000000;
	sineTable[10'd289] = 26'b01100100001000100111110101;
	sineTable[10'd290] = 26'b11111111111110111111111111;
	sineTable[10'd291] = 26'b10011011110110100111110101;
	sineTable[10'd292] = 26'b10000000000011111111111111;
	sineTable[10'd293] = 26'b10011011110110100111110101;
	sineTable[10'd294] = 26'b11111111111110111111111111;
	sineTable[10'd295] = 26'b01100100001000100111110101;
	sineTable[10'd296] = 26'b01111111111110000000000000;
	sineTable[10'd297] = 26'b01100100001000100111110101;
	sineTable[10'd298] = 26'b11111111111110111111111111;
	sineTable[10'd299] = 26'b10011011110110100111110101;
	sineTable[10'd300] = 26'b10000000000011111111111111;
	sineTable[10'd301] = 26'b10011011110111011000001010;
	sineTable[10'd302] = 26'b00000000000001000000000001;
	sineTable[10'd303] = 26'b01100100001001011000001010;
	sineTable[10'd304] = 26'b01111111111110000000000000;
	sineTable[10'd305] = 26'b01100100001000100111110101;
	sineTable[10'd306] = 26'b11111111111110111111111111;
	sineTable[10'd307] = 26'b10011011110110100111110101;
	sineTable[10'd308] = 26'b10000000000011111111111111;
	sineTable[10'd309] = 26'b10011011110110100111110101;
	sineTable[10'd310] = 26'b11111111111110111111111111;
	sineTable[10'd311] = 26'b01100100001000100111110101;
	sineTable[10'd312] = 26'b01111111111110000000000000;
	sineTable[10'd313] = 26'b01100100001001011000001010;
	sineTable[10'd314] = 26'b00000000000001000000000001;
	sineTable[10'd315] = 26'b10011011110111011000001010;
	sineTable[10'd316] = 26'b10000000000011111111111111;
	sineTable[10'd317] = 26'b10011011110110100111110101;
	sineTable[10'd318] = 26'b11111111111110111111111111;
	sineTable[10'd319] = 26'b01100100001000100111110101;
	sineTable[10'd320] = 26'b01111111111110000000000000;
	sineTable[10'd321] = 26'b01100100001001011000001010;
	sineTable[10'd322] = 26'b00000000000001000000000001;
	sineTable[10'd323] = 26'b10011011110111011000001010;
	sineTable[10'd324] = 26'b10000000000011111111111111;
	sineTable[10'd325] = 26'b10011011110110100111110101;
	sineTable[10'd326] = 26'b11111111111110111111111111;
	sineTable[10'd327] = 26'b01100100001000100111110101;
	sineTable[10'd328] = 26'b01111111111110000000000000;
	sineTable[10'd329] = 26'b01100100001000100111110101;
	sineTable[10'd330] = 26'b11111111111110111111111111;
	sineTable[10'd331] = 26'b10011011110110100111110101;
	sineTable[10'd332] = 26'b10000000000011111111111111;
	sineTable[10'd333] = 26'b10011011110110100111110101;
	sineTable[10'd334] = 26'b11111111111110111111111111;
	sineTable[10'd335] = 26'b01100100001000100111110101;
	sineTable[10'd336] = 26'b01111111111110000000000000;
	sineTable[10'd337] = 26'b01100100001000100111110101;
	sineTable[10'd338] = 26'b11111111111110111111111111;
	sineTable[10'd339] = 26'b10011011110110100111110101;
	sineTable[10'd340] = 26'b10000000000011111111111111;
	sineTable[10'd341] = 26'b10011011110111011000001010;
	sineTable[10'd342] = 26'b00000000000001000000000001;
	sineTable[10'd343] = 26'b01100100001001011000001010;
	sineTable[10'd344] = 26'b01111111111110000000000000;
	sineTable[10'd345] = 26'b01100100001000100111110101;
	sineTable[10'd346] = 26'b11111111111110111111111111;
	sineTable[10'd347] = 26'b10011011110110100111110101;
	sineTable[10'd348] = 26'b10000000000011111111111111;
	sineTable[10'd349] = 26'b10011011110110100111110101;
	sineTable[10'd350] = 26'b11111111111110111111111111;
	sineTable[10'd351] = 26'b01100100001000100111110101;
	sineTable[10'd352] = 26'b01111111111110000000000000;
	sineTable[10'd353] = 26'b01100100001000100111110101;
	sineTable[10'd354] = 26'b11111111111110111111111111;
	sineTable[10'd355] = 26'b10011011110110100111110101;
	sineTable[10'd356] = 26'b10000000000011111111111111;
	sineTable[10'd357] = 26'b10011011110110100111110101;
	sineTable[10'd358] = 26'b11111111111110111111111111;
	sineTable[10'd359] = 26'b01100100001000100111110101;
	sineTable[10'd360] = 26'b01111111111110000000000000;
	sineTable[10'd361] = 26'b01100100001001011000001010;
	sineTable[10'd362] = 26'b00000000000001000000000001;
	sineTable[10'd363] = 26'b10011011110111011000001010;
	sineTable[10'd364] = 26'b10000000000011111111111111;
	sineTable[10'd365] = 26'b10011011110110100111110101;
	sineTable[10'd366] = 26'b11111111111110111111111111;
	sineTable[10'd367] = 26'b01100100001000100111110101;
	sineTable[10'd368] = 26'b01111111111110000000000000;
	sineTable[10'd369] = 26'b01100100001001011000001010;
	sineTable[10'd370] = 26'b00000000000001000000000001;
	sineTable[10'd371] = 26'b10011011110111011000001010;
	sineTable[10'd372] = 26'b10000000000011111111111111;
	sineTable[10'd373] = 26'b10011011110111011000001010;
	sineTable[10'd374] = 26'b00000000000001000000000001;
	sineTable[10'd375] = 26'b01100100001001011000001010;
	sineTable[10'd376] = 26'b01111111111110000000000000;
	sineTable[10'd377] = 26'b01100100001000100111110101;
	sineTable[10'd378] = 26'b11111111111110111111111111;
	sineTable[10'd379] = 26'b10011011110110100111110101;
	sineTable[10'd380] = 26'b10000000000011111111111111;
	sineTable[10'd381] = 26'b10011011110111011000001010;
	sineTable[10'd382] = 26'b00000000000001000000000001;
	sineTable[10'd383] = 26'b01100100001001011000001010;
	sineTable[10'd384] = 26'b01111111111110000000000000;
	sineTable[10'd385] = 26'b01100100001001011000001010;
	sineTable[10'd386] = 26'b00000000000001000000000001;
	sineTable[10'd387] = 26'b10011011110111011000001010;
	sineTable[10'd388] = 26'b10000000000011111111111111;
	sineTable[10'd389] = 26'b10011011110110100111110101;
	sineTable[10'd390] = 26'b11111111111110111111111111;
	sineTable[10'd391] = 26'b01100100001000100111110101;
	sineTable[10'd392] = 26'b01111111111110000000000000;
	sineTable[10'd393] = 26'b01100100001000100111110101;
	sineTable[10'd394] = 26'b11111111111110111111111111;
	sineTable[10'd395] = 26'b10011011110110100111110101;
	sineTable[10'd396] = 26'b10000000000011111111111111;
	sineTable[10'd397] = 26'b10011011110111011000001010;
	sineTable[10'd398] = 26'b00000000000001000000000001;
	sineTable[10'd399] = 26'b01100100001001011000001010;
	sineTable[10'd400] = 26'b01111111111110000000000000;
	sineTable[10'd401] = 26'b01100100001000100111110101;
	sineTable[10'd402] = 26'b11111111111110111111111111;
	sineTable[10'd403] = 26'b10011011110110100111110101;
	sineTable[10'd404] = 26'b10000000000011111111111111;
	sineTable[10'd405] = 26'b10011011110110100111110101;
	sineTable[10'd406] = 26'b11111111111110111111111111;
	sineTable[10'd407] = 26'b01100100001000100111110101;
	sineTable[10'd408] = 26'b01111111111110000000000000;
	sineTable[10'd409] = 26'b01100100001000100111110101;
	sineTable[10'd410] = 26'b11111111111110111111111111;
	sineTable[10'd411] = 26'b10011011110110100111110101;
	sineTable[10'd412] = 26'b10000000000011111111111111;
	sineTable[10'd413] = 26'b10011011110110100111110101;
	sineTable[10'd414] = 26'b11111111111110111111111111;
	sineTable[10'd415] = 26'b01100100001000100111110101;
	sineTable[10'd416] = 26'b01111111111110000000000000;
	sineTable[10'd417] = 26'b01100100001001011000001010;
	sineTable[10'd418] = 26'b00000000000001000000000001;
	sineTable[10'd419] = 26'b10011011110111011000001010;
	sineTable[10'd420] = 26'b10000000000011111111111111;
	sineTable[10'd421] = 26'b10011011110111011000001010;
	sineTable[10'd422] = 26'b00000000000001000000000001;
	sineTable[10'd423] = 26'b01100100001001011000001010;
	sineTable[10'd424] = 26'b01111111111110000000000000;
	sineTable[10'd425] = 26'b01100100001001011000001010;
	sineTable[10'd426] = 26'b00000000000001000000000001;
	sineTable[10'd427] = 26'b10011011110111011000001010;
	sineTable[10'd428] = 26'b10000000000011111111111111;
	sineTable[10'd429] = 26'b10011011110110100111110101;
	sineTable[10'd430] = 26'b11111111111110111111111111;
	sineTable[10'd431] = 26'b01100100001000100111110101;
	sineTable[10'd432] = 26'b01111111111110000000000000;
	sineTable[10'd433] = 26'b01100100001000100111110101;
	sineTable[10'd434] = 26'b11111111111110111111111111;
	sineTable[10'd435] = 26'b10011011110110100111110101;
	sineTable[10'd436] = 26'b10000000000011111111111111;
	sineTable[10'd437] = 26'b10011011110110100111110101;
	sineTable[10'd438] = 26'b11111111111110111111111111;
	sineTable[10'd439] = 26'b01100100001000100111110101;
	sineTable[10'd440] = 26'b01111111111110000000000000;
	sineTable[10'd441] = 26'b01100100001000100111110101;
	sineTable[10'd442] = 26'b11111111111110111111111111;
	sineTable[10'd443] = 26'b10011011110110100111110101;
	sineTable[10'd444] = 26'b10000000000011111111111111;
	sineTable[10'd445] = 26'b10011011110110100111110101;
	sineTable[10'd446] = 26'b11111111111110111111111111;
	sineTable[10'd447] = 26'b01100100001000100111110101;
	sineTable[10'd448] = 26'b01111111111110000000000000;
	sineTable[10'd449] = 26'b01100100001001011000001010;
	sineTable[10'd450] = 26'b00000000000001000000000001;
	sineTable[10'd451] = 26'b10011011110111011000001010;
	sineTable[10'd452] = 26'b10000000000011111111111111;
	sineTable[10'd453] = 26'b10011011110110100111110101;
	sineTable[10'd454] = 26'b11111111111110111111111111;
	sineTable[10'd455] = 26'b01100100001000100111110101;
	sineTable[10'd456] = 26'b01111111111110000000000000;
	sineTable[10'd457] = 26'b01100100001000100111110101;
	sineTable[10'd458] = 26'b11111111111110111111111111;
	sineTable[10'd459] = 26'b10011011110110100111110101;
	sineTable[10'd460] = 26'b10000000000011111111111111;
	sineTable[10'd461] = 26'b10011011110111011000001010;
	sineTable[10'd462] = 26'b00000000000001000000000001;
	sineTable[10'd463] = 26'b01100100001001011000001010;
	sineTable[10'd464] = 26'b01111111111110000000000000;
	sineTable[10'd465] = 26'b01100100001000100111110101;
	sineTable[10'd466] = 26'b11111111111110111111111111;
	sineTable[10'd467] = 26'b10011011110110100111110101;
	sineTable[10'd468] = 26'b10000000000011111111111111;
	sineTable[10'd469] = 26'b10011011110111011000001010;
	sineTable[10'd470] = 26'b00000000000001000000000001;
	sineTable[10'd471] = 26'b01100100001001011000001010;
	sineTable[10'd472] = 26'b01111111111110000000000000;
	sineTable[10'd473] = 26'b01100100001001011000001010;
	sineTable[10'd474] = 26'b00000000000001000000000001;
	sineTable[10'd475] = 26'b10011011110111011000001010;
	sineTable[10'd476] = 26'b10000000000011111111111111;
	sineTable[10'd477] = 26'b10011011110111011000001010;
	sineTable[10'd478] = 26'b00000000000001000000000001;
	sineTable[10'd479] = 26'b01100100001001011000001010;
	sineTable[10'd480] = 26'b01111111111110000000000000;
	sineTable[10'd481] = 26'b01100100001001011000001010;
	sineTable[10'd482] = 26'b00000000000001000000000001;
	sineTable[10'd483] = 26'b10011011110111011000001010;
	sineTable[10'd484] = 26'b10000000000011111111111111;
	sineTable[10'd485] = 26'b10011011110111011000001010;
	sineTable[10'd486] = 26'b00000000000001000000000001;
	sineTable[10'd487] = 26'b01100100001001011000001010;
	sineTable[10'd488] = 26'b01111111111110000000000000;
	sineTable[10'd489] = 26'b01100100001000100111110101;
	sineTable[10'd490] = 26'b11111111111110111111111111;
	sineTable[10'd491] = 26'b10011011110110100111110101;
	sineTable[10'd492] = 26'b10000000000011111111111111;
	sineTable[10'd493] = 26'b10011011110111011000001010;
	sineTable[10'd494] = 26'b00000000000001000000000001;
	sineTable[10'd495] = 26'b01100100001001011000001010;
	sineTable[10'd496] = 26'b01111111111110000000000000;
	sineTable[10'd497] = 26'b01100100001000100111110101;
	sineTable[10'd498] = 26'b11111111111110111111111111;
	sineTable[10'd499] = 26'b10011011110110100111110101;
	sineTable[10'd500] = 26'b10000000000011111111111111;
	sineTable[10'd501] = 26'b10011011110110100111110101;
	sineTable[10'd502] = 26'b11111111111110111111111111;
	sineTable[10'd503] = 26'b01100100001000100111110101;
	sineTable[10'd504] = 26'b01111111111110000000000000;
	sineTable[10'd505] = 26'b01100100001001011000001010;
	sineTable[10'd506] = 26'b00000000000001000000000001;
	sineTable[10'd507] = 26'b10011011110111011000001010;
	sineTable[10'd508] = 26'b10000000000011111111111111;
	sineTable[10'd509] = 26'b10011011110111011000001010;
	sineTable[10'd510] = 26'b00000000000001000000000001;
	sineTable[10'd511] = 26'b01100100001001011000001010;
	sineTable[10'd512] = 26'b01111111111110000000000000;
	sineTable[10'd513] = 26'b01100100001001011000001010;
	sineTable[10'd514] = 26'b00000000000001000000000001;
	sineTable[10'd515] = 26'b10011011110111011000001010;
	sineTable[10'd516] = 26'b10000000000011111111111111;
	sineTable[10'd517] = 26'b10011011110111011000001010;
	sineTable[10'd518] = 26'b00000000000001000000000001;
	sineTable[10'd519] = 26'b01100100001001011000001010;
	sineTable[10'd520] = 26'b01111111111110000000000000;
	sineTable[10'd521] = 26'b01100100001001011000001010;
	sineTable[10'd522] = 26'b00000000000001000000000001;
	sineTable[10'd523] = 26'b10011011110111011000001010;
	sineTable[10'd524] = 26'b10000000000011111111111111;
	sineTable[10'd525] = 26'b10011011110110100111110101;
	sineTable[10'd526] = 26'b11111111111110111111111111;
	sineTable[10'd527] = 26'b01100100001000100111110101;
	sineTable[10'd528] = 26'b01111111111110000000000000;
	sineTable[10'd529] = 26'b01100100001000100111110101;
	sineTable[10'd530] = 26'b11111111111110111111111111;
	sineTable[10'd531] = 26'b10011011110110100111110101;
	sineTable[10'd532] = 26'b10000000000011111111111111;
	sineTable[10'd533] = 26'b10011011110111011000001010;
	sineTable[10'd534] = 26'b00000000000001000000000001;
	sineTable[10'd535] = 26'b01100100001001011000001010;
	sineTable[10'd536] = 26'b01111111111110000000000000;
	sineTable[10'd537] = 26'b01100100001001011000001010;
	sineTable[10'd538] = 26'b00000000000001000000000001;
	sineTable[10'd539] = 26'b10011011110111011000001010;
	sineTable[10'd540] = 26'b10000000000011111111111111;
	sineTable[10'd541] = 26'b10011011110111011000001010;
	sineTable[10'd542] = 26'b00000000000001000000000001;
	sineTable[10'd543] = 26'b01100100001001011000001010;
	sineTable[10'd544] = 26'b01111111111110000000000000;
	sineTable[10'd545] = 26'b01100100001000100111110101;
	sineTable[10'd546] = 26'b11111111111110111111111111;
	sineTable[10'd547] = 26'b10011011110110100111110101;
	sineTable[10'd548] = 26'b10000000000011111111111111;
	sineTable[10'd549] = 26'b10011011110110100111110101;
	sineTable[10'd550] = 26'b11111111111110111111111111;
	sineTable[10'd551] = 26'b01100100001000100111110101;
	sineTable[10'd552] = 26'b01111111111110000000000000;
	sineTable[10'd553] = 26'b01100100001001011000001010;
	sineTable[10'd554] = 26'b00000000000001000000000001;
	sineTable[10'd555] = 26'b10011011110111011000001010;
	sineTable[10'd556] = 26'b10000000000011111111111111;
	sineTable[10'd557] = 26'b10011011110110100111110101;
	sineTable[10'd558] = 26'b11111111111110111111111111;
	sineTable[10'd559] = 26'b01100100001000100111110101;
	sineTable[10'd560] = 26'b01111111111110000000000000;
	sineTable[10'd561] = 26'b01100100001000100111110101;
	sineTable[10'd562] = 26'b11111111111110111111111111;
	sineTable[10'd563] = 26'b10011011110110100111110101;
	sineTable[10'd564] = 26'b10000000000011111111111111;
	sineTable[10'd565] = 26'b10011011110111011000001010;
	sineTable[10'd566] = 26'b00000000000001000000000001;
	sineTable[10'd567] = 26'b01100100001001011000001010;
	sineTable[10'd568] = 26'b01111111111110000000000000;
	sineTable[10'd569] = 26'b01100100001001011000001010;
	sineTable[10'd570] = 26'b00000000000001000000000001;
	sineTable[10'd571] = 26'b10011011110111011000001010;
	sineTable[10'd572] = 26'b10000000000011111111111111;
	sineTable[10'd573] = 26'b10011011110110100111110101;
	sineTable[10'd574] = 26'b11111111111110111111111111;
	sineTable[10'd575] = 26'b01100100001000100111110101;
	sineTable[10'd576] = 26'b01111111111110000000000000;
	sineTable[10'd577] = 26'b01100100001001011000001010;
	sineTable[10'd578] = 26'b00000000000001000000000001;
	sineTable[10'd579] = 26'b10011011110111011000001010;
	sineTable[10'd580] = 26'b10000000000011111111111111;
	sineTable[10'd581] = 26'b10011011110110100111110101;
	sineTable[10'd582] = 26'b11111111111110111111111111;
	sineTable[10'd583] = 26'b01100100001000100111110101;
	sineTable[10'd584] = 26'b01111111111110000000000000;
	sineTable[10'd585] = 26'b01100100001000100111110101;
	sineTable[10'd586] = 26'b11111111111110111111111111;
	sineTable[10'd587] = 26'b10011011110110100111110101;
	sineTable[10'd588] = 26'b10000000000011111111111111;
	sineTable[10'd589] = 26'b10011011110111011000001010;
	sineTable[10'd590] = 26'b00000000000001000000000001;
	sineTable[10'd591] = 26'b01100100001001011000001010;
	sineTable[10'd592] = 26'b01111111111110000000000000;
	sineTable[10'd593] = 26'b01100100001000100111110101;
	sineTable[10'd594] = 26'b11111111111110111111111111;
	sineTable[10'd595] = 26'b10011011110110100111110101;
	sineTable[10'd596] = 26'b10000000000011111111111111;
	sineTable[10'd597] = 26'b10011011110110100111110101;
	sineTable[10'd598] = 26'b11111111111110111111111111;
	sineTable[10'd599] = 26'b01100100001000100111110101;
	sineTable[10'd600] = 26'b01111111111110000000000000;
	sineTable[10'd601] = 26'b01100100001001011000001010;
	sineTable[10'd602] = 26'b00000000000001000000000001;
	sineTable[10'd603] = 26'b10011011110111011000001010;
	sineTable[10'd604] = 26'b10000000000011111111111111;
	sineTable[10'd605] = 26'b10011011110111011000001010;
	sineTable[10'd606] = 26'b00000000000001000000000001;
	sineTable[10'd607] = 26'b01100100001001011000001010;
	sineTable[10'd608] = 26'b01111111111110000000000000;
	sineTable[10'd609] = 26'b01100100001001011000001010;
	sineTable[10'd610] = 26'b00000000000001000000000001;
	sineTable[10'd611] = 26'b10011011110111011000001010;
	sineTable[10'd612] = 26'b10000000000011111111111111;
	sineTable[10'd613] = 26'b10011011110110100111110101;
	sineTable[10'd614] = 26'b11111111111110111111111111;
	sineTable[10'd615] = 26'b01100100001000100111110101;
	sineTable[10'd616] = 26'b01111111111110000000000000;
	sineTable[10'd617] = 26'b01100100001000100111110101;
	sineTable[10'd618] = 26'b11111111111110111111111111;
	sineTable[10'd619] = 26'b10011011110110100111110101;
	sineTable[10'd620] = 26'b10000000000011111111111111;
	sineTable[10'd621] = 26'b10011011110111011000001010;
	sineTable[10'd622] = 26'b00000000000001000000000001;
	sineTable[10'd623] = 26'b01100100001001011000001010;
	sineTable[10'd624] = 26'b01111111111110000000000000;
	sineTable[10'd625] = 26'b01100100001001011000001010;
	sineTable[10'd626] = 26'b00000000000001000000000001;
	sineTable[10'd627] = 26'b10011011110111011000001010;
	sineTable[10'd628] = 26'b10000000000011111111111111;
	sineTable[10'd629] = 26'b10011011110110100111110101;
	sineTable[10'd630] = 26'b11111111111110111111111111;
	sineTable[10'd631] = 26'b01100100001000100111110101;
	sineTable[10'd632] = 26'b01111111111110000000000000;
	sineTable[10'd633] = 26'b01100100001001011000001010;
	sineTable[10'd634] = 26'b00000000000001000000000001;
	sineTable[10'd635] = 26'b10011011110111011000001010;
	sineTable[10'd636] = 26'b10000000000011111111111111;
	sineTable[10'd637] = 26'b10011011110110100111110101;
	sineTable[10'd638] = 26'b11111111111110111111111111;
	sineTable[10'd639] = 26'b01100100001000100111110101;
	sineTable[10'd640] = 26'b01111111111110000000000000;
	sineTable[10'd641] = 26'b01100100001000100111110101;
	sineTable[10'd642] = 26'b11111111111110111111111111;
	sineTable[10'd643] = 26'b10011011110110100111110101;
	sineTable[10'd644] = 26'b10000000000011111111111111;
	sineTable[10'd645] = 26'b10011011110111011000001010;
	sineTable[10'd646] = 26'b00000000000001000000000001;
	sineTable[10'd647] = 26'b01100100001001011000001010;
	sineTable[10'd648] = 26'b01111111111110000000000000;
	sineTable[10'd649] = 26'b01100100001001011000001010;
	sineTable[10'd650] = 26'b00000000000001000000000001;
	sineTable[10'd651] = 26'b10011011110111011000001010;
	sineTable[10'd652] = 26'b10000000000011111111111111;
	sineTable[10'd653] = 26'b10011011110111011000001010;
	sineTable[10'd654] = 26'b00000000000001000000000001;
	sineTable[10'd655] = 26'b01100100001001011000001010;
	sineTable[10'd656] = 26'b01111111111110000000000000;
	sineTable[10'd657] = 26'b01100100001000100111110101;
	sineTable[10'd658] = 26'b11111111111110111111111111;
	sineTable[10'd659] = 26'b10011011110110100111110101;
	sineTable[10'd660] = 26'b10000000000011111111111111;
	sineTable[10'd661] = 26'b10011011110110100111110101;
	sineTable[10'd662] = 26'b11111111111110111111111111;
	sineTable[10'd663] = 26'b01100100001000100111110101;
	sineTable[10'd664] = 26'b01111111111110000000000000;
	sineTable[10'd665] = 26'b01100100001001011000001010;
	sineTable[10'd666] = 26'b00000000000001000000000001;
	sineTable[10'd667] = 26'b10011011110111011000001010;
	sineTable[10'd668] = 26'b10000000000011111111111111;
	sineTable[10'd669] = 26'b10011011110111011000001010;
	sineTable[10'd670] = 26'b00000000000001000000000001;
	sineTable[10'd671] = 26'b01100100001001011000001010;
	sineTable[10'd672] = 26'b01111111111110000000000000;
	sineTable[10'd673] = 26'b01100100001001011000001010;
	sineTable[10'd674] = 26'b00000000000001000000000001;
	sineTable[10'd675] = 26'b10011011110111011000001010;
	sineTable[10'd676] = 26'b10000000000011111111111111;
	sineTable[10'd677] = 26'b10011011110110100111110101;
	sineTable[10'd678] = 26'b11111111111110111111111111;
	sineTable[10'd679] = 26'b01100100001000100111110101;
	sineTable[10'd680] = 26'b01111111111110000000000000;
	sineTable[10'd681] = 26'b01100100001000100111110101;
	sineTable[10'd682] = 26'b11111111111110111111111111;
	sineTable[10'd683] = 26'b10011011110110100111110101;
	sineTable[10'd684] = 26'b10000000000011111111111111;
	sineTable[10'd685] = 26'b10011011110110100111110101;
	sineTable[10'd686] = 26'b11111111111110111111111111;
	sineTable[10'd687] = 26'b01100100001000100111110101;
	sineTable[10'd688] = 26'b01111111111110000000000000;
	sineTable[10'd689] = 26'b01100100001000100111110101;
	sineTable[10'd690] = 26'b11111111111110111111111111;
	sineTable[10'd691] = 26'b10011011110110100111110101;
	sineTable[10'd692] = 26'b10000000000011111111111111;
	sineTable[10'd693] = 26'b10011011110110100111110101;
	sineTable[10'd694] = 26'b11111111111110111111111111;
	sineTable[10'd695] = 26'b01100100001000100111110101;
	sineTable[10'd696] = 26'b01111111111110000000000000;
	sineTable[10'd697] = 26'b01100100001000100111110101;
	sineTable[10'd698] = 26'b11111111111110111111111111;
	sineTable[10'd699] = 26'b10011011110110100111110101;
	sineTable[10'd700] = 26'b10000000000011111111111111;
	sineTable[10'd701] = 26'b10011011110111011000001010;
	sineTable[10'd702] = 26'b00000000000001000000000001;
	sineTable[10'd703] = 26'b01100100001001011000001010;
	sineTable[10'd704] = 26'b01111111111110000000000000;
	sineTable[10'd705] = 26'b01100100001000100111110101;
	sineTable[10'd706] = 26'b11111111111110111111111111;
	sineTable[10'd707] = 26'b10011011110110100111110101;
	sineTable[10'd708] = 26'b10000000000011111111111111;
	sineTable[10'd709] = 26'b10011011110111011000001010;
	sineTable[10'd710] = 26'b00000000000001000000000001;
	sineTable[10'd711] = 26'b01100100001001011000001010;
	sineTable[10'd712] = 26'b01111111111110000000000000;
	sineTable[10'd713] = 26'b01100100001000100111110101;
	sineTable[10'd714] = 26'b11111111111110111111111111;
	sineTable[10'd715] = 26'b10011011110110100111110101;
	sineTable[10'd716] = 26'b10000000000011111111111111;
	sineTable[10'd717] = 26'b10011011110110100111110101;
	sineTable[10'd718] = 26'b11111111111110111111111111;
	sineTable[10'd719] = 26'b01100100001000100111110101;
	sineTable[10'd720] = 26'b01111111111110000000000000;
	sineTable[10'd721] = 26'b01100100001001011000001010;
	sineTable[10'd722] = 26'b00000000000001000000000001;
	sineTable[10'd723] = 26'b10011011110111011000001010;
	sineTable[10'd724] = 26'b10000000000011111111111111;
	sineTable[10'd725] = 26'b10011011110110100111110101;
	sineTable[10'd726] = 26'b11111111111110111111111111;
	sineTable[10'd727] = 26'b01100100001000100111110101;
	sineTable[10'd728] = 26'b01111111111110000000000000;
	sineTable[10'd729] = 26'b01100100001001011000001010;
	sineTable[10'd730] = 26'b00000000000001000000000001;
	sineTable[10'd731] = 26'b10011011110111011000001010;
	sineTable[10'd732] = 26'b10000000000011111111111111;
	sineTable[10'd733] = 26'b10011011110110100111110101;
	sineTable[10'd734] = 26'b11111111111110111111111111;
	sineTable[10'd735] = 26'b01100100001000100111110101;
	sineTable[10'd736] = 26'b01111111111110000000000000;
	sineTable[10'd737] = 26'b01100100001001011000001010;
	sineTable[10'd738] = 26'b00000000000001000000000001;
	sineTable[10'd739] = 26'b10011011110111011000001010;
	sineTable[10'd740] = 26'b10000000000011111111111111;
	sineTable[10'd741] = 26'b10011011110111011000001010;
	sineTable[10'd742] = 26'b00000000000001000000000001;
	sineTable[10'd743] = 26'b01100100001001011000001010;
	sineTable[10'd744] = 26'b01111111111110000000000000;
	sineTable[10'd745] = 26'b01100100001000100111110101;
	sineTable[10'd746] = 26'b11111111111110111111111111;
	sineTable[10'd747] = 26'b10011011110110100111110101;
	sineTable[10'd748] = 26'b10000000000011111111111111;
	sineTable[10'd749] = 26'b10011011110110100111110101;
	sineTable[10'd750] = 26'b11111111111110111111111111;
	sineTable[10'd751] = 26'b01100100001000100111110101;
	sineTable[10'd752] = 26'b01111111111110000000000000;
	sineTable[10'd753] = 26'b01100100001000100111110101;
	sineTable[10'd754] = 26'b11111111111110111111111111;
	sineTable[10'd755] = 26'b10011011110110100111110101;
	sineTable[10'd756] = 26'b10000000000011111111111111;
	sineTable[10'd757] = 26'b10011011110111011000001010;
	sineTable[10'd758] = 26'b00000000000001000000000001;
	sineTable[10'd759] = 26'b01100100001001011000001010;
	sineTable[10'd760] = 26'b01111111111110000000000000;
	sineTable[10'd761] = 26'b01100100001001011000001010;
	sineTable[10'd762] = 26'b00000000000001000000000001;
	sineTable[10'd763] = 26'b10011011110111011000001010;
	sineTable[10'd764] = 26'b10000000000011111111111111;
	sineTable[10'd765] = 26'b10011011110111011000001010;
	sineTable[10'd766] = 26'b00000000000001000000000001;
	sineTable[10'd767] = 26'b01100100001001011000001010;
	sineTable[10'd768] = 26'b01111111111110000000000000;
	sineTable[10'd769] = 26'b01100100001001011000001010;
	sineTable[10'd770] = 26'b00000000000001000000000001;
	sineTable[10'd771] = 26'b10011011110111011000001010;
	sineTable[10'd772] = 26'b10000000000011111111111111;
	sineTable[10'd773] = 26'b10011011110110100111110101;
	sineTable[10'd774] = 26'b11111111111110111111111111;
	sineTable[10'd775] = 26'b01100100001000100111110101;
	sineTable[10'd776] = 26'b01111111111110000000000000;
	sineTable[10'd777] = 26'b01100100001000100111110101;
	sineTable[10'd778] = 26'b11111111111110111111111111;
	sineTable[10'd779] = 26'b10011011110110100111110101;
	sineTable[10'd780] = 26'b10000000000011111111111111;
	sineTable[10'd781] = 26'b10011011110111011000001010;
	sineTable[10'd782] = 26'b00000000000001000000000001;
	sineTable[10'd783] = 26'b01100100001001011000001010;
	sineTable[10'd784] = 26'b01111111111110000000000000;
	sineTable[10'd785] = 26'b01100100001000100111110101;
	sineTable[10'd786] = 26'b11111111111110111111111111;
	sineTable[10'd787] = 26'b10011011110110100111110101;
	sineTable[10'd788] = 26'b10000000000011111111111111;
	sineTable[10'd789] = 26'b10011011110111011000001010;
	sineTable[10'd790] = 26'b00000000000001000000000001;
	sineTable[10'd791] = 26'b01100100001001011000001010;
	sineTable[10'd792] = 26'b01111111111110000000000000;
	sineTable[10'd793] = 26'b01100100001000100111110101;
	sineTable[10'd794] = 26'b11111111111110111111111111;
	sineTable[10'd795] = 26'b10011011110110100111110101;
	sineTable[10'd796] = 26'b10000000000011111111111111;
	sineTable[10'd797] = 26'b10011011110110100111110101;
	sineTable[10'd798] = 26'b11111111111110111111111111;
	sineTable[10'd799] = 26'b01100100001000100111110101;
	sineTable[10'd800] = 26'b01111111111110000000000000;
	sineTable[10'd801] = 26'b01100100001000100111110101;
	sineTable[10'd802] = 26'b11111111111110111111111111;
	sineTable[10'd803] = 26'b10011011110110100111110101;
	sineTable[10'd804] = 26'b10000000000011111111111111;
	sineTable[10'd805] = 26'b10011011110111011000001010;
	sineTable[10'd806] = 26'b00000000000001000000000001;
	sineTable[10'd807] = 26'b01100100001001011000001010;
	sineTable[10'd808] = 26'b01111111111110000000000000;
	sineTable[10'd809] = 26'b01100100001001011000001010;
	sineTable[10'd810] = 26'b00000000000001000000000001;
	sineTable[10'd811] = 26'b10011011110111011000001010;
	sineTable[10'd812] = 26'b10000000000011111111111111;
	sineTable[10'd813] = 26'b10011011110110100111110101;
	sineTable[10'd814] = 26'b11111111111110111111111111;
	sineTable[10'd815] = 26'b01100100001000100111110101;
	sineTable[10'd816] = 26'b01111111111110000000000000;
	sineTable[10'd817] = 26'b01100100001001011000001010;
	sineTable[10'd818] = 26'b00000000000001000000000001;
	sineTable[10'd819] = 26'b10011011110111011000001010;
	sineTable[10'd820] = 26'b10000000000011111111111111;
	sineTable[10'd821] = 26'b10011011110111011000001010;
	sineTable[10'd822] = 26'b00000000000001000000000001;
	sineTable[10'd823] = 26'b01100100001001011000001010;
	sineTable[10'd824] = 26'b01111111111110000000000000;
	sineTable[10'd825] = 26'b01100100001000100111110101;
	sineTable[10'd826] = 26'b11111111111110111111111111;
	sineTable[10'd827] = 26'b10011011110110100111110101;
	sineTable[10'd828] = 26'b10000000000011111111111111;
	sineTable[10'd829] = 26'b10011011110110100111110101;
	sineTable[10'd830] = 26'b11111111111110111111111111;
	sineTable[10'd831] = 26'b01100100001000100111110101;
	sineTable[10'd832] = 26'b01111111111110000000000000;
	sineTable[10'd833] = 26'b01100100001000100111110101;
	sineTable[10'd834] = 26'b11111111111110111111111111;
	sineTable[10'd835] = 26'b10011011110110100111110101;
	sineTable[10'd836] = 26'b10000000000011111111111111;
	sineTable[10'd837] = 26'b10011011110111011000001010;
	sineTable[10'd838] = 26'b00000000000001000000000001;
	sineTable[10'd839] = 26'b01100100001001011000001010;
	sineTable[10'd840] = 26'b01111111111110000000000000;
	sineTable[10'd841] = 26'b01100100001000100111110101;
	sineTable[10'd842] = 26'b11111111111110111111111111;
	sineTable[10'd843] = 26'b10011011110110100111110101;
	sineTable[10'd844] = 26'b10000000000011111111111111;
	sineTable[10'd845] = 26'b10011011110110100111110101;
	sineTable[10'd846] = 26'b11111111111110111111111111;
	sineTable[10'd847] = 26'b01100100001000100111110101;
	sineTable[10'd848] = 26'b01111111111110000000000000;
	sineTable[10'd849] = 26'b01100100001000100111110101;
	sineTable[10'd850] = 26'b11111111111110111111111111;
	sineTable[10'd851] = 26'b10011011110110100111110101;
	sineTable[10'd852] = 26'b10000000000011111111111111;
	sineTable[10'd853] = 26'b10011011110110100111110101;
	sineTable[10'd854] = 26'b11111111111110111111111111;
	sineTable[10'd855] = 26'b01100100001000100111110101;
	sineTable[10'd856] = 26'b01111111111110000000000000;
	sineTable[10'd857] = 26'b01100100001000100111110101;
	sineTable[10'd858] = 26'b11111111111110111111111111;
	sineTable[10'd859] = 26'b10011011110110100111110101;
	sineTable[10'd860] = 26'b10000000000011111111111111;
	sineTable[10'd861] = 26'b10011011110110100111110101;
	sineTable[10'd862] = 26'b11111111111110111111111111;
	sineTable[10'd863] = 26'b01100100001000100111110101;
	sineTable[10'd864] = 26'b01111111111110000000000000;
	sineTable[10'd865] = 26'b01100100001000100111110101;
	sineTable[10'd866] = 26'b11111111111110111111111111;
	sineTable[10'd867] = 26'b10011011110110100111110101;
	sineTable[10'd868] = 26'b10000000000011111111111111;
	sineTable[10'd869] = 26'b10011011110110100111110101;
	sineTable[10'd870] = 26'b11111111111110111111111111;
	sineTable[10'd871] = 26'b01100100001000100111110101;
	sineTable[10'd872] = 26'b01111111111110000000000000;
	sineTable[10'd873] = 26'b01100100001000100111110101;
	sineTable[10'd874] = 26'b11111111111110111111111111;
	sineTable[10'd875] = 26'b10011011110110100111110101;
	sineTable[10'd876] = 26'b10000000000011111111111111;
	sineTable[10'd877] = 26'b10011011110111011000001010;
	sineTable[10'd878] = 26'b00000000000001000000000001;
	sineTable[10'd879] = 26'b01100100001001011000001010;
	sineTable[10'd880] = 26'b01111111111110000000000000;
	sineTable[10'd881] = 26'b01100100001000100111110101;
	sineTable[10'd882] = 26'b11111111111110111111111111;
	sineTable[10'd883] = 26'b10011011110110100111110101;
	sineTable[10'd884] = 26'b10000000000011111111111111;
	sineTable[10'd885] = 26'b10011011110110100111110101;
	sineTable[10'd886] = 26'b11111111111110111111111111;
	sineTable[10'd887] = 26'b01100100001000100111110101;
	sineTable[10'd888] = 26'b01111111111110000000000000;
	sineTable[10'd889] = 26'b01100100001001011000001010;
	sineTable[10'd890] = 26'b00000000000001000000000001;
	sineTable[10'd891] = 26'b10011011110111011000001010;
	sineTable[10'd892] = 26'b10000000000011111111111111;
	sineTable[10'd893] = 26'b10011011110110100111110101;
	sineTable[10'd894] = 26'b11111111111110111111111111;
	sineTable[10'd895] = 26'b01100100001000100111110101;
	sineTable[10'd896] = 26'b01111111111110000000000000;
	sineTable[10'd897] = 26'b01100100001001011000001010;
	sineTable[10'd898] = 26'b00000000000001000000000001;
	sineTable[10'd899] = 26'b10011011110111011000001010;
	sineTable[10'd900] = 26'b10000000000011111111111111;
	sineTable[10'd901] = 26'b10011011110111011000001010;
	sineTable[10'd902] = 26'b00000000000001000000000001;
	sineTable[10'd903] = 26'b01100100001001011000001010;
	sineTable[10'd904] = 26'b01111111111110000000000000;
	sineTable[10'd905] = 26'b01100100001001011000001010;
	sineTable[10'd906] = 26'b00000000000001000000000001;
	sineTable[10'd907] = 26'b10011011110111011000001010;
	sineTable[10'd908] = 26'b10000000000011111111111111;
	sineTable[10'd909] = 26'b10011011110110100111110101;
	sineTable[10'd910] = 26'b11111111111110111111111111;
	sineTable[10'd911] = 26'b01100100001000100111110101;
	sineTable[10'd912] = 26'b01111111111110000000000000;
	sineTable[10'd913] = 26'b01100100001001011000001010;
	sineTable[10'd914] = 26'b00000000000001000000000001;
	sineTable[10'd915] = 26'b10011011110111011000001010;
	sineTable[10'd916] = 26'b10000000000011111111111111;
	sineTable[10'd917] = 26'b10011011110110100111110101;
	sineTable[10'd918] = 26'b11111111111110111111111111;
	sineTable[10'd919] = 26'b01100100001000100111110101;
	sineTable[10'd920] = 26'b01111111111110000000000000;
	sineTable[10'd921] = 26'b01100100001000100111110101;
	sineTable[10'd922] = 26'b11111111111110111111111111;
	sineTable[10'd923] = 26'b10011011110110100111110101;
	sineTable[10'd924] = 26'b10000000000011111111111111;
	sineTable[10'd925] = 26'b10011011110110100111110101;
	sineTable[10'd926] = 26'b11111111111110111111111111;
	sineTable[10'd927] = 26'b01100100001000100111110101;
	sineTable[10'd928] = 26'b01111111111110000000000000;
	sineTable[10'd929] = 26'b01100100001000100111110101;
	sineTable[10'd930] = 26'b11111111111110111111111111;
	sineTable[10'd931] = 26'b10011011110110100111110101;
	sineTable[10'd932] = 26'b10000000000011111111111111;
	sineTable[10'd933] = 26'b10011011110110100111110101;
	sineTable[10'd934] = 26'b11111111111110111111111111;
	sineTable[10'd935] = 26'b01100100001000100111110101;
	sineTable[10'd936] = 26'b01111111111110000000000000;
	sineTable[10'd937] = 26'b01100100001000100111110101;
	sineTable[10'd938] = 26'b11111111111110111111111111;
	sineTable[10'd939] = 26'b10011011110110100111110101;
	sineTable[10'd940] = 26'b10000000000011111111111111;
	sineTable[10'd941] = 26'b10011011110110100111110101;
	sineTable[10'd942] = 26'b11111111111110111111111111;
	sineTable[10'd943] = 26'b01100100001000100111110101;
	sineTable[10'd944] = 26'b01111111111110000000000000;
	sineTable[10'd945] = 26'b01100100001001011000001010;
	sineTable[10'd946] = 26'b00000000000001000000000001;
	sineTable[10'd947] = 26'b10011011110111011000001010;
	sineTable[10'd948] = 26'b10000000000011111111111111;
	sineTable[10'd949] = 26'b10011011110110100111110101;
	sineTable[10'd950] = 26'b11111111111110111111111111;
	sineTable[10'd951] = 26'b01100100001000100111110101;
	sineTable[10'd952] = 26'b01111111111110000000000000;
	sineTable[10'd953] = 26'b01100100001000100111110101;
	sineTable[10'd954] = 26'b11111111111110111111111111;
	sineTable[10'd955] = 26'b10011011110110100111110101;
	sineTable[10'd956] = 26'b10000000000011111111111111;
	sineTable[10'd957] = 26'b10011011110111011000001010;
	sineTable[10'd958] = 26'b00000000000001000000000001;
	sineTable[10'd959] = 26'b01100100001001011000001010;
	sineTable[10'd960] = 26'b01111111111110000000000000;
	sineTable[10'd961] = 26'b01100100001000100111110101;
	sineTable[10'd962] = 26'b11111111111110111111111111;
	sineTable[10'd963] = 26'b10011011110110100111110101;
	sineTable[10'd964] = 26'b10000000000011111111111111;
	sineTable[10'd965] = 26'b10011011110110100111110101;
	sineTable[10'd966] = 26'b11111111111110111111111111;
	sineTable[10'd967] = 26'b01100100001000100111110101;
	sineTable[10'd968] = 26'b01111111111110000000000000;
	sineTable[10'd969] = 26'b01100100001001011000001010;
	sineTable[10'd970] = 26'b00000000000001000000000001;
	sineTable[10'd971] = 26'b10011011110111011000001010;
	sineTable[10'd972] = 26'b10000000000011111111111111;
	sineTable[10'd973] = 26'b10011011110111011000001010;
	sineTable[10'd974] = 26'b00000000000001000000000001;
	sineTable[10'd975] = 26'b01100100001001011000001010;
	sineTable[10'd976] = 26'b01111111111110000000000000;
	sineTable[10'd977] = 26'b01100100001000100111110101;
	sineTable[10'd978] = 26'b11111111111110111111111111;
	sineTable[10'd979] = 26'b10011011110110100111110101;
	sineTable[10'd980] = 26'b10000000000011111111111111;
	sineTable[10'd981] = 26'b10011011110111011000001010;
	sineTable[10'd982] = 26'b00000000000001000000000001;
	sineTable[10'd983] = 26'b01100100001001011000001010;
	sineTable[10'd984] = 26'b01111111111110000000000000;
	sineTable[10'd985] = 26'b01100100001001011000001010;
	sineTable[10'd986] = 26'b00000000000001000000000001;
	sineTable[10'd987] = 26'b10011011110111011000001010;
	sineTable[10'd988] = 26'b10000000000011111111111111;
	sineTable[10'd989] = 26'b10011011110111011000001010;
	sineTable[10'd990] = 26'b00000000000001000000000001;
	sineTable[10'd991] = 26'b01100100001001011000001010;
	sineTable[10'd992] = 26'b01111111111110000000000000;
	sineTable[10'd993] = 26'b01100100001001011000001010;
	sineTable[10'd994] = 26'b00000000000001000000000001;
	sineTable[10'd995] = 26'b10011011110111011000001010;
	sineTable[10'd996] = 26'b10000000000011111111111111;
	sineTable[10'd997] = 26'b10011011110111011000001010;
	sineTable[10'd998] = 26'b00000000000001000000000001;
	sineTable[10'd999] = 26'b01100100001001011000001010;
	sineTable[10'd1000] = 26'b01111111111110000000000000;
	sineTable[10'd1001] = 26'b01100100001001011000001010;
	sineTable[10'd1002] = 26'b00000000000001000000000001;
	sineTable[10'd1003] = 26'b10011011110111011000001010;
	sineTable[10'd1004] = 26'b10000000000011111111111111;
	sineTable[10'd1005] = 26'b10011011110111011000001010;
	sineTable[10'd1006] = 26'b00000000000001000000000001;
	sineTable[10'd1007] = 26'b01100100001001011000001010;
	sineTable[10'd1008] = 26'b01111111111110000000000000;
	sineTable[10'd1009] = 26'b01100100001001011000001010;
	sineTable[10'd1010] = 26'b00000000000001000000000001;
	sineTable[10'd1011] = 26'b10011011110111011000001010;
	sineTable[10'd1012] = 26'b10000000000011111111111111;
	sineTable[10'd1013] = 26'b10011011110110100111110101;
	sineTable[10'd1014] = 26'b11111111111110111111111111;
	sineTable[10'd1015] = 26'b01100100001000100111110101;
	sineTable[10'd1016] = 26'b01111111111110000000000000;
	sineTable[10'd1017] = 26'b01100100001000100111110101;
	sineTable[10'd1018] = 26'b11111111111110111111111111;
	sineTable[10'd1019] = 26'b10011011110110100111110101;
	sineTable[10'd1020] = 26'b10000000000011111111111111;
	sineTable[10'd1021] = 26'b10011011110110100111110101;
	sineTable[10'd1022] = 26'b11111111111110111111111111;
	sineTable[10'd1023] = 26'b01100100001000100111110101;
end
endmodule
