/* Verilog model created from schematic test.sch -- May 09, 2019 15:49 */

module test;




endmodule // test
