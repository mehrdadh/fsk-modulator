/* Verilog model created from schematic test.sch -- May 14, 2019 16:13 */

module test;




endmodule // test
